44	4
shingles	yghg	zgzg	CeBe	CeCe	mgCe	Beme	aame	Reme	yeye	mexe	xeTg	ReRe	yexe	o5xe	Tgme	xeme	mgng	meCe	mezg	Q5xe	aaCg	Tgxe	yeCe	yeme	yeCg	ye	meye	ogye	aaTg	Q5Re	xeye	xexe	aaxe	me	mera	yeRe	Bezg	Tgye	xeDa	zg	Cexe	aaDa	meme	Daye
1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	1	0	0	0	1	0	0	0	1	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
2	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	2	0	0	0	0	0	1	0	1	0	2	0	0	0	0	0	0	2	0	1	0	0	1	0	0	0	0	1	0
0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	2	1	0	0	1	0	1	0	0	1	0	1	0	1	0	0	1	0	0	0	0	0
5	0	0	0	0	0	0	0	1	1	0	1	1	2	1	1	0	0	0	0	1	0	0	0	0	0	0	1	0	0	1	4	0	0	0	0	0	0	1	0	0	0	1	1	1
3	0	1	2	1	0	1	1	0	0	1	0	0	0	0	0	1	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	1	0	0	0	0	2	0	0	1	1	0	0	0
4	1	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0
